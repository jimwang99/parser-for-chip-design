**********************************************************************

.GLOBAL DVDD DVSS 
.SUBCKT CLK_GEN WENA RENA CLK CLK_ WCK RCK SEN

X2 CLK_D1 CLK_1      INV_D1
X3 RE_P CLK_D1 CLK_1 NOR2
X4 CLK_1 CLK         BUF_1
X5 WCK  WE_I WE_P    NOR2
X6 NET2 RE_I RE_P    NAND2
X7 WE_I WENA           INV
X9 WE_P CLK_1 CLK_D1 NAND2
X10 RE_I RENA CLK CLK_ FF

X8A RCK  NET2         INV_D2
X8B NET2C  RCK         INV
X8C SEN  NET2C         INV

.ENDS


.SUBCKT INV Z A LP=0.18u WP=2.40u LN=0.18u WN=1.20u
MI1 Z A DVDD DVDD TP W=WP L=LP
MI2 Z A DVSS DVSS TN W=WN L=LN
.ENDS


.SUBCKT INV_D1 Z A 
MI1 N1 A  DVDD DVDD TP W=1.20u L=0.18u
MI2 N1 A  DVSS DVSS TN W=0.60u L=0.18u
ML1 DVDD N1 DVDD DVDD TP W=5.0u L=0.36u
ML2 DVSS N1 DVSS DVSS TN W=5.0u L=0.36u
MI3 N2 N1 DVDD DVDD TP W=0.30u L=0.20u
MI4 N2 N1 DVSS DVSS TN W=0.20u L=0.20u
ML3 DVDD N2 DVDD DVDD TP W=5.0u L=0.36u
ML4 DVSS N2 DVSS DVSS TN W=5.0u L=0.36u
MI5 N3 N2 DVDD DVDD TP W=0.30u L=0.20u
MI6 N3 N2 DVSS DVSS TN W=0.20u L=0.20u
ML5 DVDD N3 DVDD DVDD TP W=5.0u L=0.36u
ML6 DVSS N3 DVSS DVSS TN W=5.0u L=0.36u
MI7 N4 N3 DVDD DVDD TP W=0.30u L=0.20u
MI8 N4 N3 DVSS DVSS TN W=0.20u L=0.20u
ML7 DVDD N4 DVDD DVDD TP W=5.0u L=0.36u
ML8 DVSS N4 DVSS DVSS TN W=5.0u L=0.36u
MI9 Z  N4 DVDD DVDD TP W=2.40u L=0.18u
MIA Z  N4 DVSS DVSS TN W=1.20u L=0.18u
.ENDS


.SUBCKT INV_D2 Z A 
MI1 N1 A  DVDD DVDD TP W=1.20u L=0.18u
MI2 N1 A  DVSS DVSS TN W=0.60u L=0.18u
ML1 DVDD N1 DVDD DVDD TP W=2.0u L=0.36u
ML2 DVSS N1 DVSS DVSS TN W=1.0u L=0.36u
MI3 N2 N1 DVDD DVDD TP W=0.30u L=0.20u
MI4 N2 N1 DVSS DVSS TN W=0.20u L=0.20u
ML3 DVDD N2 DVDD DVDD TP W=5.0u L=0.36u
ML4 DVSS N2 DVSS DVSS TN W=5.0u L=0.36u
MI5 N3 N2 DVDD DVDD TP W=0.30u L=0.20u
MI6 N3 N2 DVSS DVSS TN W=0.20u L=0.20u
ML5 DVDD N3 DVDD DVDD TP W=5.0u L=0.36u
ML6 DVSS N3 DVSS DVSS TN W=5.0u L=0.36u
MI7 N4 N3 DVDD DVDD TP W=0.30u L=0.20u
MI8 N4 N3 DVSS DVSS TN W=0.20u L=0.20u
ML7 DVDD N4 DVDD DVDD TP W=5.0u L=0.36u
ML8 DVSS N4 DVSS DVSS TN W=5.0u L=0.36u
MI9 Z  N4 DVDD DVDD TP W=2.40u L=0.18u
MIA Z  N4 DVSS DVSS TN W=1.20u L=0.18u
.ENDS



.SUBCKT BUF_1 Z A LN=0.18u LP=0.18u WN=1.20u WP=0.60u
MP1 NET1 A DVDD DVDD TP W=WP L=LP
MN1 NET1 A DVSS DVSS TN W=WN L=LN
MP2 Z NET1 DVDD DVDD TP W=WP L=LP
MN2 Z NET1 DVSS DVSS TN W=WN L=LN
.ENDS


.SUBCKT DEC A_2_ A_1_ A_0_ WCK RCK CLK CLK_ 
+ WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_

X1 AD_2_ A_2_ CLK CLK_ FF
X2 AD_1_ A_1_ CLK CLK_ FF
X3 AD_0_ A_0_ CLK CLK_ FF
X4 XAD_2_ AD_2_ INV
X5 XAD_1_ AD_1_ INV
X6 XAD_0_ AD_0_ INV
X7 WCK_ WCK INV
X8 RCK_ RCK INV
XD7 W_7_ AD_2_  AD_1_  AD_0_  NAND3
XD6 W_6_ AD_2_  AD_1_  XAD_0_ NAND3
XD5 W_5_ AD_2_  XAD_1_ AD_0_  NAND3
XD4 W_4_ AD_2_  XAD_1_ XAD_0_ NAND3
XD3 W_3_ XAD_2_ AD_1_  AD_0_  NAND3
XD2 W_2_ XAD_2_ AD_1_  XAD_0_ NAND3
XD1 W_1_ XAD_2_ XAD_1_ AD_0_  NAND3
XD0 W_0_ XAD_2_ XAD_1_ XAD_0_ NAND3
XE7 WWL_7_ W_7_ WCK_ NOR2
XE6 WWL_6_ W_6_ WCK_ NOR2
XE5 WWL_5_ W_5_ WCK_ NOR2
XE4 WWL_4_ W_4_ WCK_ NOR2
XE3 WWL_3_ W_3_ WCK_ NOR2
XE2 WWL_2_ W_2_ WCK_ NOR2
XE1 WWL_1_ W_1_ WCK_ NOR2
XE0 WWL_0_ W_0_ WCK_ NOR2
XF7 RWL_7_ W_7_ RCK_ RNOR22
XF6 RWL_6_ W_6_ RCK_ RNOR22
XF5 RWL_5_ W_5_ RCK_ RNOR22
XF4 RWL_4_ W_4_ RCK_ RNOR22
XF3 RWL_3_ W_3_ RCK_ RNOR22
XF2 RWL_2_ W_2_ RCK_ RNOR22
XF1 RWL_1_ W_1_ RCK_ RNOR22
XF0 RWL_0_ W_0_ RCK_ RNOR22
.ENDS


.SUBCKT NOR2 Z A B 
+ LPA=0.18u LNA=0.18u LPB=0.18u LNB=0.18u
+ WPA=4.80u WNA=1.20u WPB=4.80u WNB=1.20u
MI1 NET1 A DVDD DVDD TP W=WPA L=LPA
MI2 Z B NET1    DVDD TP W=WPB L=LPB
MI3 Z A DVSS    DVSS TN W=WNA L=LNA
MI4 Z B DVSS    DVSS TN W=WNB L=LNB
.ENDS

.SUBCKT RNOR22 Z A B 
+ LPA=0.18u LNA=0.18u LPB=0.18u LNB=0.18u
+ WPA=4.80u WNA=1.20u WPB=4.80u WNB=1.20u
MI1 NET1 A DVDD DVDD TP W=WPA L=LPA
MI2 Z B NET1    DVDD TP W=WPB L=LPB
MI3 Z A DVSS    DVSS TN W=WNA L=LNA
MI4 Z B DVSS    DVSS TN W=WNB L=LNB
.ENDS

.SUBCKT WNOR22 Z A B
+ LPA=0.18u LNA=0.18u LPB=0.18u LNB=0.18u
+ WPA=2.40u WNA=2.40u WPB=2.40u WNB=2.40u
MP1 Z A DVDD    DVDD TP W=WPA L=LPA 
MP2 Z B DVDD    DVDD TP W=WPB L=LPB 
MN1 Z A NET1    DVSS TN W=WNA L=LNA 
MN2 NET1 B DVSS DVSS TN W=WNB L=LNB 
.ENDS

.SUBCKT NAND2 Z A B
+ LPA=0.18u LNA=0.18u LPB=0.18u LNB=0.18u
+ WPA=2.40u WNA=2.40u WPB=2.40u WNB=2.40u
MP1 Z A DVDD    DVDD TP W=WPA L=LPA 
MP2 Z B DVDD    DVDD TP W=WPB L=LPB 
MN1 Z A NET1    DVSS TN W=WNA L=LNA 
MN2 NET1 B DVSS DVSS TN W=WNB L=LNB 
.ENDS

.SUBCKT NAND3 Z A B C
+ LPA=0.18u LNA=0.18u LPB=0.18u LNB=0.18u LPC=0.18u LNC=0.18u
+ WPA=2.40u WNA=3.60u WPB=2.40u WNB=3.60u WPC=2.40u WNC=3.60u
MP1 Z A DVDD     DVDD TP W=WPA L=LPA
MP2 Z B DVDD     DVDD TP W=WPB L=LPB
MP3 Z C DVDD     DVDD TP W=WPC L=LPC
MN1 Z A NET1     DVSS TN W=WNA L=LNA
MN2 NET1 B NET2  DVSS TN W=WNB L=LNB
MN3 NET2 C DVSS  DVSS TN W=WNC L=LNC
.ENDS

.SUBCKT LAT Q D CLK

X1 CLK_ CLK INV

MP1 S CLK_ D DVDD TP L=0.18u W=2.4u
MN1 S CLK  D DVSS TN L=0.18u W=2.4u
MP2 S XQ DVDD DVDD TP L=0.18u W=1.2u
MN2 S XQ DVSS DVSS TN L=0.18u W=0.6u
MP3 XQ S DVDD DVDD TP L=0.18u W=1.2u
MN3 XQ S DVSS DVSS TN L=0.18u W=1.2u
MP4 Q XQ DVDD DVDD TP L=0.18u W=2.4u
MN4 Q XQ DVSS DVSS TN L=0.18u W=1.2u


.ENDS

.SUBCKT FF Q D CLK CLK_

X1 Q1 D  CLK_ LAT
X2 Q  Q1 CLK  LAT

.ENDS


.SUBCKT MEM WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_7_ WBL_6_ WBL_5_ WBL_4_ WBL_3_ WBL_2_ WBL_1_ WBL_0_ 
+ XWBL_7_ XWBL_6_ XWBL_5_ XWBL_4_ XWBL_3_ XWBL_2_ XWBL_1_ XWBL_0_ 
+ RBL_7_ RBL_6_ RBL_5_ RBL_4_ RBL_3_ RBL_2_ RBL_1_ RBL_0_ 
+ XRBL_7_ XRBL_6_ XRBL_5_ XRBL_4_ XRBL_3_ XRBL_2_ XRBL_1_ XRBL_0_ 

XBANK0 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_1_ XWBL_1_ RBL_1_ XRBL_1_ 
+ WBL_0_ XWBL_0_ RBL_0_ XRBL_0_ MEMBANK

XBANK1 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_3_ XWBL_3_ RBL_3_ XRBL_3_ 
+ WBL_2_ XWBL_2_ RBL_2_ XRBL_2_ MEMBANK

XBANK2 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_5_ XWBL_5_ RBL_5_ XRBL_5_ 
+ WBL_4_ XWBL_4_ RBL_4_ XRBL_4_ MEMBANK

XBANK3 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_7_ XWBL_7_ RBL_7_ XRBL_7_ 
+ WBL_6_ XWBL_6_ RBL_6_ XRBL_6_ MEMBANK

.ENDS


.SUBCKT MEMBANK WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_1_ XWBL_1_ RBL_1_ XRBL_1_ 
+ WBL_0_ XWBL_0_ RBL_0_ XRBL_0_

X0 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_0_ XWBL_0_ RBL_0_ XRBL_0_ MEMCOL
X1 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_  
+ WBL_1_ XWBL_1_ RBL_1_ XRBL_1_ MEMCOL

.ENDS


.SUBCKT MEMCOL WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL XWBL RBL XRBL

X7 WWL_7_ RWL_7_ WBL XWBL RBL XRBL MEMCELL
X6 WWL_6_ RWL_6_ WBL XWBL RBL XRBL MEMCELL
X5 WWL_5_ RWL_5_ WBL XWBL RBL XRBL MEMCELL
X4 WWL_4_ RWL_4_ WBL XWBL RBL XRBL MEMCELL
X3 WWL_3_ RWL_3_ WBL XWBL RBL XRBL MEMCELL
X2 WWL_2_ RWL_2_ WBL XWBL RBL XRBL MEMCELL
X1 WWL_1_ RWL_1_ WBL XWBL RBL XRBL MEMCELL
X0 WWL_0_ RWL_0_ WBL XWBL RBL XRBL MEMCELL

.ENDS


.SUBCKT MEMCELL WWL RWL WBL XWBL RBL XRBL 

MN1 S  WWL WBL  DVSS TN L=0.18u W=0.50u
MN2 XS WWL XWBL DVSS TN L=0.18u W=0.50u
MN3 RBL  RWL S  DVSS TN L=0.18u W=0.50u 
MN4 XRBL RWL XS DVSS TN L=0.18u W=0.50u 
MP1 XS S DVDD    DVDD TP L=0.18u W=0.50u
MP2 S XS DVDD    DVDD TP L=0.18u W=0.50u
MN5 XS S DVSS    DVSS TN L=0.18u W=1.00u
MN6 S XS DVSS    DVSS TN L=0.18u W=1.00u

.ENDS


.SUBCKT IO DI_7_ DI_6_ DI_5_ DI_4_ DI_3_ DI_2_ DI_1_ DI_0_
+ DOUT_7_ DOUT_6_ DOUT_5_ DOUT_4_ DOUT_3_ DOUT_2_ DOUT_1_ DOUT_0_ 
+ WCK RCK SEN OE XCLR
+ WBL_7_ WBL_6_ WBL_5_ WBL_4_ WBL_3_ WBL_2_ WBL_1_ WBL_0_ 
+ XWBL_7_ XWBL_6_ XWBL_5_ XWBL_4_ XWBL_3_ XWBL_2_ XWBL_1_ XWBL_0_ 
+ RBL_7_ RBL_6_ RBL_5_ RBL_4_ RBL_3_ RBL_2_ RBL_1_ RBL_0_ 
+ XRBL_7_ XRBL_6_ XRBL_5_ XRBL_4_ XRBL_3_ XRBL_2_ XRBL_1_ XRBL_0_
+ RAW_RENA RAW_OE

XW0 DI_0_ WCK WBL_0_ XWBL_0_ WDRV
XW1 DI_1_ WCK WBL_1_ XWBL_1_ WDRV
XW2 DI_2_ WCK WBL_2_ XWBL_2_ WDRV
XW3 DI_3_ WCK WBL_3_ XWBL_3_ WDRV
XW4 DI_4_ WCK WBL_4_ XWBL_4_ WDRV
XW5 DI_5_ WCK WBL_5_ XWBL_5_ WDRV
XW6 DI_6_ WCK WBL_6_ XWBL_6_ WDRV
XW7 DI_7_ WCK WBL_7_ XWBL_7_ WDRV

XR0 XDO0 SEN RBL_0_ XRBL_0_ SENSEAMP
XR1 XDO1 SEN RBL_1_ XRBL_1_ SENSEAMP
XR2 XDO2 SEN RBL_2_ XRBL_2_ SENSEAMP
XR3 XDO3 SEN RBL_3_ XRBL_3_ SENSEAMP
XR4 XDO4 SEN RBL_4_ XRBL_4_ SENSEAMP
XR5 XDO5 SEN RBL_5_ XRBL_5_ SENSEAMP
XR6 XDO6 SEN RBL_6_ XRBL_6_ SENSEAMP
XR7 XDO7 SEN RBL_7_ XRBL_7_ SENSEAMP

XOUT0 XDO0 OE XCLR DOUT_0_ RAW_RENA RAW_OE OUTBUF
XOUT1 XDO1 OE XCLR DOUT_1_ RAW_RENA RAW_OE OUTBUF
XOUT2 XDO2 OE XCLR DOUT_2_ RAW_RENA RAW_OE OUTBUF
XOUT3 XDO3 OE XCLR DOUT_3_ RAW_RENA RAW_OE OUTBUF
XOUT4 XDO4 OE XCLR DOUT_4_ RAW_RENA RAW_OE OUTBUF
XOUT5 XDO5 OE XCLR DOUT_5_ RAW_RENA RAW_OE OUTBUF
XOUT6 XDO6 OE XCLR DOUT_6_ RAW_RENA RAW_OE OUTBUF
XOUT7 XDO7 OE XCLR DOUT_7_ RAW_RENA RAW_OE OUTBUF

.ENDS

.SUBCKT WDRV DI WCK BL XBL

X1 XDI DI INV
MP1 BL WCK DVDD   DVDD TP L=0.18u W=1.2u
MP2 BL WCK XBL   DVDD TP L=0.18u W=0.8u
MP3 XBL WCK DVDD  DVDD TP L=0.18u W=1.2u
MP4 BL XBL DVDD   DVDD TP L=0.18u W=1.5u
MP5 XBL BL DVDD   DVDD TP L=0.18u W=1.5u
MN1 XBL DI NET1  DVSS TN L=0.18u W=2.4u
MN2 BL XDI NET1  DVSS TN L=0.18u W=2.4u
MN3 NET1 WCK DVSS DVSS TN L=0.18u W=1.2u

.ENDS


.SUBCKT SENSEAMP XDO SEN BL XBL

MPP1 BL SEN DVDD    DVDD TP L=0.18u W=0.8u
MPP2 XBL SEN DVDD    DVDD TP L=0.18u W=0.8u


MP1 DOUT SEN DVDD    DVDD TP L=0.18u W=0.8u
MP2 DOUT SEN XDOUT    DVDD TP L=0.18u W=0.8u
MP3 XDOUT SEN DVDD   DVDD TP L=0.18u W=0.8u
MP6 DOUT XDOUT DVDD    DVDD TP L=0.18u W=1.5u
MP7 XDOUT DOUT DVDD    DVDD TP L=0.18u W=1.5u

MN10 DOUT XBL N1 DVSS TN L=0.18u W=1.5u
MN11 XDOUT BL N1 DVSS TN L=0.18u W=1.5u
MN12 N1  SEN DVSS  DVSS TN L=0.18u W=1.5u

MN13 XDO SEN XDOUT DVSS TN L=0.18u W=3.0u

.ENDS

.SUBCKT OUTBUF XDO OE XCLR DOUT RAW_RENA RAW_OE

X1 XOE OE INV LP=0.18u WP=2.40u LN=0.18u WN=1.20u

MP1 NS XOE XDO DVDD TP L=0.18u W=4.0u
MN1 NS OE XDO DVSS TN L=0.18u W=2.0u

MP3 NS DOUTI DVDD DVDD TP L=0.18u W=0.60u
MN3 NS DOUTI DVSS DVSS TN L=0.18u W=0.30u

MP4 DOUTI NS DVDD DVDD TP L=0.18u W=2.40u
MN4 DOUTI NS DVSS DVSS TN L=0.18u W=1.20u

MP5 NS XCLR DVDD DVDD TP L=0.18u W=0.70u

*MP6 NS OE   DVDD DVDD TP L=0.18u W=0.80u
X2 XDOUT DOUTI  RAW_RENA  RAW_OE  NAND3
X3 DOUT XDOUT INV

.ENDS


.SUBCKT RAM1R1W A<2> A<1> A<0> DI<7> DI<6> DI<5> DI<4> DI<3> DI<2> DI<1> DI<0>
+ DOUT<7> DOUT<6> DOUT<5> DOUT<4> DOUT<3> DOUT<2> DOUT<1> DOUT<0> WENA RENA OE CLR CLK

XI1 WENA RENA CLK CLK_ WCK RCK SEN CLK_GEN
XI2 A<2> A<1> A<0> WCK RCK CLK CLK_ 
+ WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ DEC
XI4 CLK_ CLK INV
XI5 WWL_7_ WWL_6_ WWL_5_ WWL_4_ WWL_3_ WWL_2_ WWL_1_ WWL_0_ 
+ RWL_7_ RWL_6_ RWL_5_ RWL_4_ RWL_3_ RWL_2_ RWL_1_ RWL_0_ 
+ WBL_7_ WBL_6_ WBL_5_ WBL_4_ WBL_3_ WBL_2_ WBL_1_ WBL_0_ 
+ XWBL_7_ XWBL_6_ XWBL_5_ XWBL_4_ XWBL_3_ XWBL_2_ XWBL_1_ XWBL_0_ 
+ RBL_7_ RBL_6_ RBL_5_ RBL_4_ RBL_3_ RBL_2_ RBL_1_ RBL_0_ 
+ XRBL_7_ XRBL_6_ XRBL_5_ XRBL_4_ XRBL_3_ XRBL_2_ XRBL_1_ XRBL_0_ 
+ MEM
XI6 D7 D6 D5 D4 D3 D2 D1 D0
+ DOUT<7> DOUT<6> DOUT<5> DOUT<4> DOUT<3> DOUT<2> DOUT<1> DOUT<0> 
+ WCK RCK SEN OE_I XCLR
+ WBL_7_ WBL_6_ WBL_5_ WBL_4_ WBL_3_ WBL_2_ WBL_1_ WBL_0_ 
+ XWBL_7_ XWBL_6_ XWBL_5_ XWBL_4_ XWBL_3_ XWBL_2_ XWBL_1_ XWBL_0_ 
+ RBL_7_ RBL_6_ RBL_5_ RBL_4_ RBL_3_ RBL_2_ RBL_1_ RBL_0_ 
+ XRBL_7_ XRBL_6_ XRBL_5_ XRBL_4_ XRBL_3_ XRBL_2_ XRBL_1_ XRBL_0_
+ RENA OE
+ IO

XDI0 D0 DI<0> CLK CLK_ FF
XDI1 D1 DI<1> CLK CLK_ FF
XDI2 D2 DI<2> CLK CLK_ FF
XDI3 D3 DI<3> CLK CLK_ FF
XDI4 D4 DI<4> CLK CLK_ FF
XDI5 D5 DI<5> CLK CLK_ FF
XDI6 D6 DI<6> CLK CLK_ FF
XDI7 D7 DI<7> CLK CLK_ FF
XOE OE_I OE CLK CLK_ FF
XCLRFF CLR_I CLR CLK CLK_ FF
XCLKD CLKD CLK_ INV
XCLRIIFF CLR_II CLR_I CLK_ CLKD FF
XCLRINV XCLR CLR_II INV

.ENDS
